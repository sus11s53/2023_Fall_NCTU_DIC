.SUBCKT Adder_1bit_FULL_ADDER VSS VDD  X Y CIN COUT SUM
XU1 VSS VDD  X Y A AND2x2_ASAP7_75t_R
XU2 VSS VDD  Y X B XOR2xp5_ASAP7_75t_R
XU3 VSS VDD  B CIN SUM XOR2xp5_ASAP7_75t_R
XU4 VSS VDD  B CIN C AND2x2_ASAP7_75t_R
XU5 VSS VDD  C CIN COUT OR2x2_ASAP7_75t_R
.ENDS


