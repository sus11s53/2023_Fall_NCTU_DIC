.SUBCKT Adder_1bit A B Output[1] Output[0]
XU1 A B Output[1] AND2x2_ASAP7_75t_R
XU2 B A Output[0] XOR2xp5_ASAP7_75t_R
.ENDS


