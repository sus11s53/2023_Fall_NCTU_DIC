//==============================================
//==============================================				
//	Author	:	Wei Lu																		
//----------------------------------------------
//												
//	File Name		:	Comparator.v					
//	Module Name		:	Comparator					
//	Release version	:	v1.0					
//----------------------------------------------										

module Comparator(
    //Input Port
	A,
	B,	
    //Output Port
	Out
    );

//---------------------------------------------------------------------
//   PORT DECLARATION
//---------------------------------------------------------------------
input[63:0]A;
input[63:0]B;
output reg Out;


//---------------------------------------------------------------------
//   Design
//---------------------------------------------------------------------
always@(*)
begin
	if(A == B)
		Out = 1'd1;
	else
		Out = 1'd0;
end



endmodule