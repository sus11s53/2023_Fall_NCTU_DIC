.SUBCKT Convolution VSS VDD  In_IFM_1[3] In_IFM_1[2] In_IFM_1[1] In_IFM_1[0] In_IFM_2[3] In_IFM_2[2] In_IFM_2[1] In_IFM_2[0] In_IFM_3[3] In_IFM_3[2] In_IFM_3[1] In_IFM_3[0] In_IFM_4[3] In_IFM_4[2] In_IFM_4[1] In_IFM_4[0] In_Weight_1[3] In_Weight_1[2] In_Weight_1[1] In_Weight_1[0] In_Weight_2[3] In_Weight_2[2] In_Weight_2[1] In_Weight_2[0] In_Weight_3[3] In_Weight_3[2] In_Weight_3[1] In_Weight_3[0] In_Weight_4[3] In_Weight_4[2] In_Weight_4[1] In_Weight_4[0] Out_OFM[9] Out_OFM[8] Out_OFM[7] Out_OFM[6] Out_OFM[5] Out_OFM[4] Out_OFM[3] Out_OFM[2] Out_OFM[1] Out_OFM[0]
XDP_OP_10J1_122_2300_U122 VSS VDD  DP_OP_10J1_122_2300_n175 DP_OP_10J1_122_2300_n181 DP_OP_10J1_122_2300_n178 DP_OP_10J1_122_2300_n153 DP_OP_10J1_122_2300_n154 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U120 VSS VDD  DP_OP_10J1_122_2300_n223 DP_OP_10J1_122_2300_n253 DP_OP_10J1_122_2300_n226 DP_OP_10J1_122_2300_n149 DP_OP_10J1_122_2300_n150 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U109 VSS VDD  DP_OP_10J1_122_2300_n219 n144 DP_OP_10J1_122_2300_n222 DP_OP_10J1_122_2300_n131 DP_OP_10J1_122_2300_n132 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U104 VSS VDD  DP_OP_10J1_122_2300_n123 DP_OP_10J1_122_2300_n151 n37 DP_OP_10J1_122_2300_n124 DP_OP_10J1_122_2300_n125 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U89 VSS VDD  DP_OP_10J1_122_2300_n137 n32 n127 DP_OP_10J1_122_2300_n101 DP_OP_10J1_122_2300_n102 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U86 VSS VDD  DP_OP_10J1_122_2300_n104 DP_OP_10J1_122_2300_n131 DP_OP_10J1_122_2300_n106 DP_OP_10J1_122_2300_n95 DP_OP_10J1_122_2300_n96 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U82 VSS VDD  DP_OP_10J1_122_2300_n99 DP_OP_10J1_122_2300_n121 n11 DP_OP_10J1_122_2300_n90 DP_OP_10J1_122_2300_n91 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U74 VSS VDD  DP_OP_10J1_122_2300_n172 DP_OP_10J1_122_2300_n241 n72 DP_OP_10J1_122_2300_n78 DP_OP_10J1_122_2300_n79 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U73 VSS VDD  DP_OP_10J1_122_2300_n196 DP_OP_10J1_122_2300_n220 n141 DP_OP_10J1_122_2300_n76 DP_OP_10J1_122_2300_n77 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U64 VSS VDD  DP_OP_10J1_122_2300_n69 DP_OP_10J1_122_2300_n72 n12 DP_OP_10J1_122_2300_n63 DP_OP_10J1_122_2300_n64 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U58 VSS VDD  DP_OP_10J1_122_2300_n192 DP_OP_10J1_122_2300_n216 DP_OP_10J1_122_2300_n80 DP_OP_10J1_122_2300_n54 DP_OP_10J1_122_2300_n55 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U56 VSS VDD  DP_OP_10J1_122_2300_n76 DP_OP_10J1_122_2300_n78 DP_OP_10J1_122_2300_n51 DP_OP_10J1_122_2300_n52 DP_OP_10J1_122_2300_n53 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U54 VSS VDD  n116 DP_OP_10J1_122_2300_n74 DP_OP_10J1_122_2300_n71 DP_OP_10J1_122_2300_n49 DP_OP_10J1_122_2300_n50 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U49 VSS VDD  DP_OP_10J1_122_2300_n52 DP_OP_10J1_122_2300_n56 n75 DP_OP_10J1_122_2300_n41 DP_OP_10J1_122_2300_n42 FAx1_ASAP7_75t_R
XDP_OP_10J1_122_2300_U48 VSS VDD  n56 DP_OP_10J1_122_2300_n49 DP_OP_10J1_122_2300_n46 DP_OP_10J1_122_2300_n38 DP_OP_10J1_122_2300_n39 FAx1_ASAP7_75t_R
XU1 VSS VDD  n251 n9 Out_OFM[7] XOR2x2_ASAP7_75t_R
XU2 VSS VDD  n249 n59 Out_OFM[5] XNOR2xp5_ASAP7_75t_R
XU3 VSS VDD  n247 n62 Out_OFM[6] XNOR2xp5_ASAP7_75t_R
XU4 VSS VDD  n85 n86 n251 XNOR2xp5_ASAP7_75t_R
XU5 VSS VDD  DP_OP_10J1_122_2300_n125 n189 n61 XNOR2xp5_ASAP7_75t_R
XU6 VSS VDD  n58 n70 n107 XOR2xp5_ASAP7_75t_R
XU7 VSS VDD  n24 n103 INVx1_ASAP7_75t_R
XU8 VSS VDD  n27 n212 INVx2_ASAP7_75t_R
XU9 VSS VDD  n123 n55 n58 XNOR2xp5_ASAP7_75t_R
XU10 VSS VDD  n82 n203 INVx2_ASAP7_75t_R
XU11 VSS VDD  DP_OP_10J1_122_2300_n125 n189 n228 XNOR2xp5_ASAP7_75t_R
XU12 VSS VDD  n28 n10 INVx2_ASAP7_75t_R
XU13 VSS VDD  n69 DP_OP_10J1_122_2300_n128 n189 XNOR2xp5_ASAP7_75t_R
XU14 VSS VDD  DP_OP_10J1_122_2300_n79 DP_OP_10J1_122_2300_n98 n178 XNOR2xp5_ASAP7_75t_R
XU15 VSS VDD  n168 n29 DP_OP_10J1_122_2300_n108 XNOR2xp5_ASAP7_75t_R
XU16 VSS VDD  n122 n142 n196 NOR2x1_ASAP7_75t_R
XU17 VSS VDD  n241 n179 n193 NOR2x1_ASAP7_75t_R
XU18 VSS VDD  n186 n25 INVx3_ASAP7_75t_R
XU19 VSS VDD  n137 n134 DP_OP_10J1_122_2300_n226 NOR2x1_ASAP7_75t_R
XU20 VSS VDD  n153 n148 n172 NOR2x1_ASAP7_75t_R
XU21 VSS VDD  n135 n138 DP_OP_10J1_122_2300_n196 NOR2xp67_ASAP7_75t_R
XU22 VSS VDD  In_IFM_4[0] In_Weight_4[1] n216 NAND2xp5_ASAP7_75t_R
XU23 VSS VDD  In_IFM_4[2] In_Weight_4[3] DP_OP_10J1_122_2300_n172 AND2x2_ASAP7_75t_R
XU24 VSS VDD  n89 n88 n177 NOR2x1_ASAP7_75t_R
XU25 VSS VDD  n18 n23 DP_OP_10J1_122_2300_n198 NOR2x1_ASAP7_75t_R
XU26 VSS VDD  In_IFM_2[0] In_Weight_2[3] DP_OP_10J1_122_2300_n204 AND2x2_ASAP7_75t_R
XU27 VSS VDD  n115 n155 DP_OP_10J1_122_2300_n205 NOR2xp67_ASAP7_75t_R
XU28 VSS VDD  DP_OP_10J1_122_2300_n153 n13 INVx1_ASAP7_75t_R
XU29 VSS VDD  n131 n236 DP_OP_10J1_122_2300_n246 NOR2xp33_ASAP7_75t_R
XU30 VSS VDD  n130 n140 DP_OP_10J1_122_2300_n245 NOR2xp33_ASAP7_75t_R
XU31 VSS VDD  n246 n1 Out_OFM[8] XNOR2x1_ASAP7_75t_R
XU32 VSS VDD  n6 n4 n5 n1 MAJIxp5_ASAP7_75t_R
XU33 VSS VDD  n13 DP_OP_10J1_122_2300_n243 DP_OP_10J1_122_2300_n246 DP_OP_10J1_122_2300_n127 MAJIxp5_ASAP7_75t_R
XU34 VSS VDD  n71 n74 DP_OP_10J1_122_2300_n128 n64 MAJIxp5_ASAP7_75t_R
XU35 VSS VDD  n2 n13 DP_OP_10J1_122_2300_n128 XOR2xp5_ASAP7_75t_R
XU36 VSS VDD  DP_OP_10J1_122_2300_n246 DP_OP_10J1_122_2300_n243 n2 XNOR2xp5_ASAP7_75t_R
XU37 VSS VDD  n3 n55 n8 XNOR2xp5_ASAP7_75t_R
XU38 VSS VDD  n64 DP_OP_10J1_122_2300_n119 n28 n55 MAJIxp5_ASAP7_75t_R
XU39 VSS VDD  n123 n3 INVx1_ASAP7_75t_R
XU40 VSS VDD  n86 n4 INVx1_ASAP7_75t_R
XU41 VSS VDD  n85 n5 INVx1_ASAP7_75t_R
XU42 VSS VDD  n34 n30 n210 n6 MAJIxp5_ASAP7_75t_R
XU43 VSS VDD  n182 n49 DP_OP_10J1_122_2300_n104 XNOR2x2_ASAP7_75t_R
XU44 VSS VDD  In_IFM_4[0] In_Weight_4[2] DP_OP_10J1_122_2300_n181 AND2x4_ASAP7_75t_R
XU45 VSS VDD  DP_OP_10J1_122_2300_n141 n226 DP_OP_10J1_122_2300_n143 n7 MAJIxp5_ASAP7_75t_R
XU46 VSS VDD  n80 n8 n35 XNOR2xp5_ASAP7_75t_R
XU47 VSS VDD  DP_OP_10J1_122_2300_n101 n178 DP_OP_10J1_122_2300_n69 XOR2x2_ASAP7_75t_R
XU48 VSS VDD  n34 n209 n210 n9 MAJIxp5_ASAP7_75t_R
XU49 VSS VDD  n111 n12 INVx3_ASAP7_75t_R
XU50 VSS VDD  DP_OP_10J1_122_2300_n96 n28 BUFx4_ASAP7_75t_R
XU51 VSS VDD  n82 n133 n14 n80 MAJx2_ASAP7_75t_R
XU52 VSS VDD  DP_OP_10J1_122_2300_n102 DP_OP_10J1_122_2300_n89 BUFx2_ASAP7_75t_R
XU53 VSS VDD  DP_OP_10J1_122_2300_n89 n11 INVx2_ASAP7_75t_R
XU54 VSS VDD  DP_OP_10J1_122_2300_n90 n111 BUFx3_ASAP7_75t_R
XU55 VSS VDD  n41 n40 n39 n37 MAJx2_ASAP7_75t_R
XU56 VSS VDD  n16 n54 n53 DP_OP_10J1_122_2300_n98 MAJx2_ASAP7_75t_R
XU57 VSS VDD  n25 n114 DP_OP_10J1_122_2300_n124 n26 MAJx2_ASAP7_75t_R
XU58 VSS VDD  n238 n237 n52 XOR2xp5_ASAP7_75t_R
XU59 VSS VDD  n214 n213 DP_OP_10J1_122_2300_n137 NOR2x1p5_ASAP7_75t_R
XU60 VSS VDD  In_IFM_4[2] In_Weight_4[1] n213 NAND2x1_ASAP7_75t_R
XU61 VSS VDD  In_Weight_1[2] In_IFM_1[0] n40 NAND2x1_ASAP7_75t_R
XU62 VSS VDD  n181 n180 n49 XOR2x1_ASAP7_75t_R
XU63 VSS VDD  DP_OP_10J1_122_2300_n120 DP_OP_10J1_122_2300_n140 DP_OP_10J1_122_2300_n122 n14 MAJIxp5_ASAP7_75t_R
XU64 VSS VDD  DP_OP_10J1_122_2300_n223 DP_OP_10J1_122_2300_n253 DP_OP_10J1_122_2300_n226 A0  n15 FAx1_ASAP7_75t_R
XU65 VSS VDD  n104 n71 INVx3_ASAP7_75t_R
XU66 VSS VDD  DP_OP_10J1_122_2300_n91 n82 BUFx4_ASAP7_75t_R
XU67 VSS VDD  n238 n237 n16 XNOR2xp5_ASAP7_75t_R
XU68 VSS VDD  In_IFM_2[0] n17 INVx8_ASAP7_75t_R
XU69 VSS VDD  In_IFM_2[2] n18 INVx8_ASAP7_75t_R
XU70 VSS VDD  In_IFM_2[0] n155 INVx8_ASAP7_75t_R
XU71 VSS VDD  In_IFM_1[2] n19 INVx8_ASAP7_75t_R
XU72 VSS VDD  In_IFM_1[2] n20 INVx8_ASAP7_75t_R
XU73 VSS VDD  DP_OP_10J1_122_2300_n40 n75 INVx4_ASAP7_75t_R
XU74 VSS VDD  DP_OP_10J1_122_2300_n54 DP_OP_10J1_122_2300_n40 BUFx5_ASAP7_75t_R
XU75 VSS VDD  DP_OP_10J1_122_2300_n38 n27 BUFx5_ASAP7_75t_R
XU76 VSS VDD  In_IFM_4[1] In_Weight_4[3] n21 AND2x2_ASAP7_75t_R
XU77 VSS VDD  DP_OP_10J1_122_2300_n39 n24 BUFx2_ASAP7_75t_R
XU78 VSS VDD  DP_OP_10J1_122_2300_n127 n186 BUFx5_ASAP7_75t_R
XU79 VSS VDD  In_Weight_2[1] n22 INVx8_ASAP7_75t_R
XU80 VSS VDD  In_Weight_2[1] n23 INVx8_ASAP7_75t_R
XU81 VSS VDD  n83 n104 BUFx4_ASAP7_75t_R
XU82 VSS VDD  n211 n33 n30 XNOR2xp5_ASAP7_75t_R
XU83 VSS VDD  In_IFM_4[1] In_Weight_4[3] n29 NAND2xp33_ASAP7_75t_R
XU84 VSS VDD  In_IFM_1[1] In_Weight_1[0] n79 AND2x2_ASAP7_75t_R
XU85 VSS VDD  n43 n44 n42 NAND2xp33_ASAP7_75t_R
XU86 VSS VDD  n172 n79 n163 XNOR2xp5_ASAP7_75t_R
XU87 VSS VDD  n185 n188 DP_OP_10J1_122_2300_n46 NAND2x1_ASAP7_75t_R
XU88 VSS VDD  In_Weight_4[0] In_IFM_4[0] n147 NAND2xp33_ASAP7_75t_R
XU89 VSS VDD  n231 n162 Out_OFM[4] XOR2xp5_ASAP7_75t_R
XU90 VSS VDD  DP_OP_10J1_122_2300_n95 n66 n31 OR2x2_ASAP7_75t_R
XU91 VSS VDD  n233 n232 DP_OP_10J1_122_2300_n56 NOR2x1_ASAP7_75t_R
XU92 VSS VDD  n207 n206 n211 XNOR2x2_ASAP7_75t_R
XU93 VSS VDD  n61 n227 n229 XOR2xp5_ASAP7_75t_R
XU94 VSS VDD  n117 n208 INVxp67_ASAP7_75t_R
XU95 VSS VDD  n160 n110 n159 XNOR2xp5_ASAP7_75t_R
XU96 VSS VDD  DP_OP_10J1_122_2300_n198 DP_OP_10J1_122_2300_n204 n176 XOR2xp5_ASAP7_75t_R
XU97 VSS VDD  In_IFM_2[3] In_Weight_2[2] n72 AND2x2_ASAP7_75t_R
XU98 VSS VDD  In_Weight_4[0] In_IFM_4[1] n215 NAND2xp5_ASAP7_75t_R
XU99 VSS VDD  In_Weight_3[3] In_IFM_3[3] n232 NAND2x1_ASAP7_75t_R
XU100 VSS VDD  In_IFM_4[3] In_Weight_4[3] n233 NAND2x1_ASAP7_75t_R
XU101 VSS VDD  In_IFM_1[1] In_Weight_1[3] n32 AND2x2_ASAP7_75t_R
XU102 VSS VDD  In_Weight_3[3] In_IFM_3[2] n234 NAND2x1_ASAP7_75t_R
XU103 VSS VDD  In_Weight_2[0] In_IFM_2[0] n191 NAND2xp5_ASAP7_75t_R
XU104 VSS VDD  In_Weight_3[0] In_IFM_3[0] n190 NAND2xp5_ASAP7_75t_R
XU105 VSS VDD  n100 n128 n158 n36 MAJIxp5_ASAP7_75t_R
XU106 VSS VDD  n55 n132 n80 n210 MAJIxp5_ASAP7_75t_R
XU107 VSS VDD  n211 n33 n209 XNOR2xp5_ASAP7_75t_R
XU108 VSS VDD  DP_OP_10J1_122_2300_n63 n208 n33 XNOR2xp5_ASAP7_75t_R
XU109 VSS VDD  n35 n36 DP_OP_10J1_122_2300_n64 n34 MAJIxp5_ASAP7_75t_R
XU110 VSS VDD  n41 n38 DP_OP_10J1_122_2300_n148 XNOR2xp5_ASAP7_75t_R
XU111 VSS VDD  n40 n39 n38 XNOR2xp5_ASAP7_75t_R
XU112 VSS VDD  In_Weight_3[1] In_IFM_3[1] n39 NAND2xp5_ASAP7_75t_R
XU113 VSS VDD  In_IFM_3[2] In_Weight_3[0] n41 NAND2xp5_ASAP7_75t_R
XU114 VSS VDD  n31 n42 n206 NAND2xp5_ASAP7_75t_R
XU115 VSS VDD  n25 n114 DP_OP_10J1_122_2300_n124 n43 MAJIxp5_ASAP7_75t_R
XU116 VSS VDD  DP_OP_10J1_122_2300_n95 n66 n44 NAND2xp5_ASAP7_75t_R
XU117 VSS VDD  n106 n45 Out_OFM[9] NAND2x1p5_ASAP7_75t_R
XU118 VSS VDD  n101 n46 n45 NAND2xp5_ASAP7_75t_R
XU119 VSS VDD  n48 n47 n46 NAND2xp5_ASAP7_75t_R
XU120 VSS VDD  n62 n209 n210 n47 MAJIxp5_ASAP7_75t_R
XU121 VSS VDD  n86 n85 n48 NAND2xp5_ASAP7_75t_R
XU122 VSS VDD  In_IFM_1[3] In_Weight_1[1] n180 AND2x2_ASAP7_75t_R
XU123 VSS VDD  In_Weight_3[1] In_IFM_3[3] n181 AND2x2_ASAP7_75t_R
XU124 VSS VDD  In_Weight_1[2] In_IFM_1[2] n182 AND2x2_ASAP7_75t_R
XU125 VSS VDD  n50 n165 n128 XOR2x2_ASAP7_75t_R
XU126 VSS VDD  DP_OP_10J1_122_2300_n119 n10 n50 XOR2xp5_ASAP7_75t_R
XU127 VSS VDD  n54 n51 DP_OP_10J1_122_2300_n99 XNOR2xp5_ASAP7_75t_R
XU128 VSS VDD  n53 n52 n51 XNOR2xp5_ASAP7_75t_R
XU129 VSS VDD  In_Weight_4[1] In_IFM_4[3] n237 NAND2xp5_ASAP7_75t_R
XU130 VSS VDD  In_Weight_4[2] In_IFM_4[2] n238 NAND2xp5_ASAP7_75t_R
XU131 VSS VDD  DP_OP_10J1_122_2300_n225 n174 DP_OP_10J1_122_2300_n249 n53 MAJIxp5_ASAP7_75t_R
XU132 VSS VDD  n93 n92 DP_OP_10J1_122_2300_n249 NOR2x1_ASAP7_75t_R
XU133 VSS VDD  n120 n125 n174 NOR2x1_ASAP7_75t_R
XU134 VSS VDD  n95 n94 DP_OP_10J1_122_2300_n225 NOR2x1_ASAP7_75t_R
XU135 VSS VDD  DP_OP_10J1_122_2300_n204 n177 DP_OP_10J1_122_2300_n198 n54 MAJIxp5_ASAP7_75t_R
XU136 VSS VDD  DP_OP_10J1_122_2300_n52 DP_OP_10J1_122_2300_n56 n75 A1  n56 FAx1_ASAP7_75t_R
XU137 VSS VDD  In_Weight_3[3] In_IFM_3[0] n144 AND2x4_ASAP7_75t_R
XU138 VSS VDD  n58 n80 n60 XOR2xp5_ASAP7_75t_R
XU139 VSS VDD  n228 n227 n7 n57 MAJIxp5_ASAP7_75t_R
XU140 VSS VDD  n158 n128 n57 n59 MAJIxp5_ASAP7_75t_R
XU141 VSS VDD  n59 n60 DP_OP_10J1_122_2300_n64 n62 MAJIxp5_ASAP7_75t_R
XU142 VSS VDD  DP_OP_10J1_122_2300_n73 DP_OP_10J1_122_2300_n105 n87 XNOR2xp5_ASAP7_75t_R
XU143 VSS VDD  In_IFM_3[1] In_Weight_3[3] n73 AND2x2_ASAP7_75t_R
XU144 VSS VDD  In_Weight_2[1] In_IFM_2[3] n169 AND2x2_ASAP7_75t_R
XU145 VSS VDD  n73 n169 n168 XNOR2xp5_ASAP7_75t_R
XU146 VSS VDD  n170 n26 n132 XNOR2xp5_ASAP7_75t_R
XU147 VSS VDD  DP_OP_10J1_122_2300_n53 n205 n187 NAND2xp33_ASAP7_75t_R
XU148 VSS VDD  In_Weight_2[2] In_IFM_2[2] n76 AND2x2_ASAP7_75t_R
XU149 VSS VDD  In_Weight_2[3] In_IFM_2[1] n77 AND2x2_ASAP7_75t_R
XU150 VSS VDD  In_Weight_3[0] In_IFM_3[1] n194 AND2x2_ASAP7_75t_R
XU151 VSS VDD  n91 DP_OP_10J1_122_2300_n136 n90 XOR2xp5_ASAP7_75t_R
XU152 VSS VDD  n87 n67 n66 XNOR2xp5_ASAP7_75t_R
XU153 VSS VDD  n149 DP_OP_10J1_122_2300_n108 n201 XNOR2xp5_ASAP7_75t_R
XU154 VSS VDD  n21 n73 n169 n63 MAJIxp5_ASAP7_75t_R
XU155 VSS VDD  n87 n67 n65 XOR2xp5_ASAP7_75t_R
XU156 VSS VDD  n71 n74 DP_OP_10J1_122_2300_n128 n165 MAJx2_ASAP7_75t_R
XU157 VSS VDD  n21 n73 n169 n67 MAJx2_ASAP7_75t_R
XU158 VSS VDD  In_Weight_2[2] n89 INVx8_ASAP7_75t_R
XU159 VSS VDD  n143 n90 n68 XOR2xp5_ASAP7_75t_R
XU160 VSS VDD  DP_OP_10J1_122_2300_n148 DP_OP_10J1_122_2300_n152 DP_OP_10J1_122_2300_n154 n69 MAJIxp5_ASAP7_75t_R
XU161 VSS VDD  n105 n102 n101 AND2x2_ASAP7_75t_R
XU162 VSS VDD  n82 n133 n14 n70 MAJIxp5_ASAP7_75t_R
XU163 VSS VDD  DP_OP_10J1_122_2300_n148 DP_OP_10J1_122_2300_n152 DP_OP_10J1_122_2300_n154 n74 MAJx2_ASAP7_75t_R
XU164 VSS VDD  DP_OP_10J1_122_2300_n48 n116 INVx4_ASAP7_75t_R
XU165 VSS VDD  n194 n196 n193 n161 MAJx2_ASAP7_75t_R
XU166 VSS VDD  DP_OP_10J1_122_2300_n223 DP_OP_10J1_122_2300_n253 DP_OP_10J1_122_2300_n226 n81 MAJx2_ASAP7_75t_R
XU167 VSS VDD  n168 n29 n114 XOR2xp5_ASAP7_75t_R
XU168 VSS VDD  n212 DP_OP_10J1_122_2300_n41 n106 OR2x2_ASAP7_75t_R
XU169 VSS VDD  DP_OP_10J1_122_2300_n50 n211 DP_OP_10J1_122_2300_n63 n78 MAJx2_ASAP7_75t_R
XU170 VSS VDD  n37 DP_OP_10J1_122_2300_n123 DP_OP_10J1_122_2300_n151 A2  n83 FAx1_ASAP7_75t_R
XU171 VSS VDD  n214 n213 DP_OP_10J1_122_2300_n123 XNOR2xp5_ASAP7_75t_R
XU172 VSS VDD  n194 n196 n193 n84 MAJIxp5_ASAP7_75t_R
XU173 VSS VDD  DP_OP_10J1_122_2300_n50 n211 DP_OP_10J1_122_2300_n63 n85 MAJIxp5_ASAP7_75t_R
XU174 VSS VDD  DP_OP_10J1_122_2300_n42 DP_OP_10J1_122_2300_n49 DP_OP_10J1_122_2300_n46 A3  n86 FAx1_ASAP7_75t_R
XU175 VSS VDD  n63 DP_OP_10J1_122_2300_n105 DP_OP_10J1_122_2300_n73 DP_OP_10J1_122_2300_n74 MAJIxp5_ASAP7_75t_R
XU176 VSS VDD  In_IFM_2[1] n88 INVx11_ASAP7_75t_R
XU177 VSS VDD  n143 DP_OP_10J1_122_2300_n136 n91 DP_OP_10J1_122_2300_n119 MAJIxp5_ASAP7_75t_R
XU178 VSS VDD  n143 n90 DP_OP_10J1_122_2300_n120 XNOR2xp5_ASAP7_75t_R
XU179 VSS VDD  n177 n176 n91 XNOR2xp5_ASAP7_75t_R
XU180 VSS VDD  In_IFM_3[1] n92 INVx8_ASAP7_75t_R
XU181 VSS VDD  In_Weight_3[2] n93 INVx8_ASAP7_75t_R
XU182 VSS VDD  In_IFM_1[1] n94 INVx8_ASAP7_75t_R
XU183 VSS VDD  In_Weight_1[2] n95 INVx8_ASAP7_75t_R
XU184 VSS VDD  DP_OP_10J1_122_2300_n249 DP_OP_10J1_122_2300_n225 n173 XOR2xp5_ASAP7_75t_R
XU185 VSS VDD  n96 n68 n227 XNOR2xp5_ASAP7_75t_R
XU186 VSS VDD  DP_OP_10J1_122_2300_n122 DP_OP_10J1_122_2300_n140 n96 XNOR2xp5_ASAP7_75t_R
XU187 VSS VDD  DP_OP_10J1_122_2300_n158 DP_OP_10J1_122_2300_n150 n97 DP_OP_10J1_122_2300_n140 MAJIxp5_ASAP7_75t_R
XU188 VSS VDD  n199 n198 n197 DP_OP_10J1_122_2300_n158 MAJIxp5_ASAP7_75t_R
XU189 VSS VDD  n161 n159 n97 XNOR2xp5_ASAP7_75t_R
XU190 VSS VDD  DP_OP_10J1_122_2300_n132 n98 DP_OP_10J1_122_2300_n122 XNOR2xp5_ASAP7_75t_R
XU191 VSS VDD  n81 DP_OP_10J1_122_2300_n130 n98 XNOR2xp5_ASAP7_75t_R
XU192 VSS VDD  DP_OP_10J1_122_2300_n148 n99 DP_OP_10J1_122_2300_n143 XOR2xp5_ASAP7_75t_R
XU193 VSS VDD  DP_OP_10J1_122_2300_n152 DP_OP_10J1_122_2300_n154 n99 XNOR2xp5_ASAP7_75t_R
XU194 VSS VDD  n227 n230 n228 n100 MAJIxp5_ASAP7_75t_R
XU195 VSS VDD  n202 n203 n158 XNOR2xp5_ASAP7_75t_R
XU196 VSS VDD  n103 n78 n102 NAND2xp5_ASAP7_75t_R
XU197 VSS VDD  n212 DP_OP_10J1_122_2300_n41 n105 NAND2xp5_ASAP7_75t_R
XU198 VSS VDD  n112 n108 n84 n143 MAJx2_ASAP7_75t_R
XU199 VSS VDD  n215 n216 n108 OR2x2_ASAP7_75t_R
XU200 VSS VDD  n227 n61 n7 n162 MAJx2_ASAP7_75t_R
XU201 VSS VDD  n84 n159 DP_OP_10J1_122_2300_n146 XNOR2xp5_ASAP7_75t_R
XU202 VSS VDD  n215 n216 n110 NOR2xp33_ASAP7_75t_R
XU203 VSS VDD  In_Weight_2[0] In_IFM_2[3] DP_OP_10J1_122_2300_n195 AND2x4_ASAP7_75t_R
XU204 VSS VDD  n172 DP_OP_10J1_122_2300_n206 n79 n112 MAJIxp5_ASAP7_75t_R
XU205 VSS VDD  In_IFM_4[0] In_Weight_4[3] n146 AND2x4_ASAP7_75t_R
XU206 VSS VDD  n158 n128 n231 XNOR2xp5_ASAP7_75t_R
XU207 VSS VDD  In_IFM_4[1] In_Weight_4[2] n113 AND2x2_ASAP7_75t_R
XU208 VSS VDD  In_IFM_4[1] In_Weight_4[2] n157 AND2x4_ASAP7_75t_R
XU209 VSS VDD  In_Weight_2[2] n115 INVx8_ASAP7_75t_R
XU210 VSS VDD  DP_OP_10J1_122_2300_n55 DP_OP_10J1_122_2300_n48 BUFx4_ASAP7_75t_R
XU211 VSS VDD  n116 DP_OP_10J1_122_2300_n74 DP_OP_10J1_122_2300_n71 A4  n117 FAx1_ASAP7_75t_R
XU212 VSS VDD  In_Weight_1[3] n118 INVx8_ASAP7_75t_R
XU213 VSS VDD  In_IFM_1[2] n119 INVx8_ASAP7_75t_R
XU214 VSS VDD  In_IFM_1[0] n120 INVx8_ASAP7_75t_R
XU215 VSS VDD  In_Weight_4[0] In_IFM_4[0] n121 AND2x2_ASAP7_75t_R
XU216 VSS VDD  In_IFM_3[0] n122 INVx8_ASAP7_75t_R
XU217 VSS VDD  n170 n26 n123 XOR2xp5_ASAP7_75t_R
XU218 VSS VDD  In_IFM_3[3] n124 INVx8_ASAP7_75t_R
XU219 VSS VDD  In_Weight_1[3] n125 INVx8_ASAP7_75t_R
XU220 VSS VDD  In_Weight_1[3] n126 INVx8_ASAP7_75t_R
XU221 VSS VDD  n146 n157 DP_OP_10J1_122_2300_n195 n127 MAJx2_ASAP7_75t_R
XU222 VSS VDD  In_IFM_1[0] n129 INVx8_ASAP7_75t_R
XU223 VSS VDD  In_IFM_3[2] n130 INVx8_ASAP7_75t_R
XU224 VSS VDD  In_IFM_3[2] n131 INVx8_ASAP7_75t_R
XU225 VSS VDD  n205 DP_OP_10J1_122_2300_n53 n185 OR2x2_ASAP7_75t_R
XU226 VSS VDD  n201 DP_OP_10J1_122_2300_n124 n133 XOR2xp5_ASAP7_75t_R
XU227 VSS VDD  In_Weight_2[0] n153 INVx8_ASAP7_75t_R
XU228 VSS VDD  In_Weight_2[0] n240 INVx8_ASAP7_75t_R
XU229 VSS VDD  In_IFM_1[1] n134 INVx8_ASAP7_75t_R
XU230 VSS VDD  In_Weight_1[0] n184 INVx8_ASAP7_75t_R
XU231 VSS VDD  In_Weight_1[0] n154 INVx8_ASAP7_75t_R
XU232 VSS VDD  In_Weight_1[0] n192 INVx8_ASAP7_75t_R
XU233 VSS VDD  In_Weight_2[3] n135 INVx8_ASAP7_75t_R
XU234 VSS VDD  In_Weight_2[3] n164 INVx8_ASAP7_75t_R
XU235 VSS VDD  In_Weight_2[1] n136 INVx8_ASAP7_75t_R
XU236 VSS VDD  In_Weight_1[1] n137 INVx8_ASAP7_75t_R
XU237 VSS VDD  In_Weight_1[1] n179 INVx8_ASAP7_75t_R
XU238 VSS VDD  In_Weight_1[1] n217 INVx8_ASAP7_75t_R
XU239 VSS VDD  In_IFM_2[2] n138 INVx8_ASAP7_75t_R
XU240 VSS VDD  In_IFM_2[2] n239 INVx8_ASAP7_75t_R
XU241 VSS VDD  In_Weight_3[2] n139 INVx8_ASAP7_75t_R
XU242 VSS VDD  In_Weight_3[2] n140 INVx8_ASAP7_75t_R
XU243 VSS VDD  In_IFM_1[3] In_Weight_1[2] n141 AND2x2_ASAP7_75t_R
XU244 VSS VDD  In_Weight_3[1] n142 INVx11_ASAP7_75t_R
XU245 VSS VDD  In_Weight_3[1] n236 INVx8_ASAP7_75t_R
XU246 VSS VDD  In_IFM_1[3] n145 INVx8_ASAP7_75t_R
XU247 VSS VDD  In_IFM_1[3] n183 INVx8_ASAP7_75t_R
XU248 VSS VDD  In_IFM_2[1] n148 INVx8_ASAP7_75t_R
XU249 VSS VDD  In_IFM_2[1] n152 INVx8_ASAP7_75t_R
XU250 VSS VDD  DP_OP_10J1_122_2300_n243 DP_OP_10J1_122_2300_n246 n13 n149 MAJIxp5_ASAP7_75t_R
XU251 VSS VDD  DP_OP_10J1_122_2300_n42 DP_OP_10J1_122_2300_n49 DP_OP_10J1_122_2300_n46 n150 MAJIxp5_ASAP7_75t_R
XU252 VSS VDD  n151 DP_OP_10J1_122_2300_n146 DP_OP_10J1_122_2300_n141 XNOR2xp5_ASAP7_75t_R
XU253 VSS VDD  n15 DP_OP_10J1_122_2300_n158 n151 XNOR2xp5_ASAP7_75t_R
XU254 VSS VDD  n172 DP_OP_10J1_122_2300_n206 n79 n160 MAJIxp5_ASAP7_75t_R
XU255 VSS VDD  n17 n22 DP_OP_10J1_122_2300_n206 NOR2x1p5_ASAP7_75t_R
XU256 VSS VDD  n146 n156 DP_OP_10J1_122_2300_n136 XNOR2xp5_ASAP7_75t_R
XU257 VSS VDD  DP_OP_10J1_122_2300_n195 n113 n156 XOR2xp5_ASAP7_75t_R
XU258 VSS VDD  DP_OP_10J1_122_2300_n206 n163 n199 XNOR2xp5_ASAP7_75t_R
XU259 VSS VDD  DP_OP_10J1_122_2300_n199 DP_OP_10J1_122_2300_n205 n167 DP_OP_10J1_122_2300_n151 MAJIxp5_ASAP7_75t_R
XU260 VSS VDD  n167 n166 DP_OP_10J1_122_2300_n152 XNOR2xp5_ASAP7_75t_R
XU261 VSS VDD  DP_OP_10J1_122_2300_n199 DP_OP_10J1_122_2300_n205 n166 XOR2xp5_ASAP7_75t_R
XU262 VSS VDD  n136 n152 n167 NOR2x1_ASAP7_75t_R
XU263 VSS VDD  DP_OP_10J1_122_2300_n95 n65 n170 XNOR2xp5_ASAP7_75t_R
XU264 VSS VDD  DP_OP_10J1_122_2300_n245 n77 n76 DP_OP_10J1_122_2300_n105 MAJIxp5_ASAP7_75t_R
XU265 VSS VDD  n77 n171 DP_OP_10J1_122_2300_n106 XNOR2xp5_ASAP7_75t_R
XU266 VSS VDD  n76 DP_OP_10J1_122_2300_n245 n171 XOR2xp5_ASAP7_75t_R
XU267 VSS VDD  DP_OP_10J1_122_2300_n141 n226 DP_OP_10J1_122_2300_n143 n230 MAJIxp5_ASAP7_75t_R
XU268 VSS VDD  n174 n173 DP_OP_10J1_122_2300_n130 XNOR2xp5_ASAP7_75t_R
XU269 VSS VDD  DP_OP_10J1_122_2300_n77 DP_OP_10J1_122_2300_n103 DP_OP_10J1_122_2300_n70 DP_OP_10J1_122_2300_n71 MAJIxp5_ASAP7_75t_R
XU270 VSS VDD  n175 DP_OP_10J1_122_2300_n77 DP_OP_10J1_122_2300_n72 XNOR2xp5_ASAP7_75t_R
XU271 VSS VDD  DP_OP_10J1_122_2300_n70 DP_OP_10J1_122_2300_n103 n175 XOR2xp5_ASAP7_75t_R
XU272 VSS VDD  DP_OP_10J1_122_2300_n132 DP_OP_10J1_122_2300_n149 DP_OP_10J1_122_2300_n130 DP_OP_10J1_122_2300_n121 MAJIxp5_ASAP7_75t_R
XU273 VSS VDD  In_Weight_3[2] n244 INVx8_ASAP7_75t_R
XU274 VSS VDD  n218 n244 DP_OP_10J1_122_2300_n241 NOR2x1_ASAP7_75t_R
XU275 VSS VDD  In_IFM_3[3] n218 INVx8_ASAP7_75t_R
XU276 VSS VDD  n20 n126 DP_OP_10J1_122_2300_n220 NOR2x1_ASAP7_75t_R
XU277 VSS VDD  n240 n239 DP_OP_10J1_122_2300_n199 NOR2x1_ASAP7_75t_R
XU278 VSS VDD  In_IFM_2[3] n243 INVx8_ASAP7_75t_R
XU279 VSS VDD  In_IFM_1[0] n241 INVx8_ASAP7_75t_R
XU280 VSS VDD  n245 n139 DP_OP_10J1_122_2300_n253 NOR2x1_ASAP7_75t_R
XU281 VSS VDD  In_IFM_3[0] n245 INVx8_ASAP7_75t_R
XU282 VSS VDD  n19 n184 DP_OP_10J1_122_2300_n223 NOR2x1_ASAP7_75t_R
XU283 VSS VDD  n119 n217 DP_OP_10J1_122_2300_n222 NOR2x1_ASAP7_75t_R
XU284 VSS VDD  n191 n190 n197 NOR2xp33_ASAP7_75t_R
XU285 VSS VDD  n216 n215 n198 XOR2xp5_ASAP7_75t_R
XU286 VSS VDD  n182 n181 n180 DP_OP_10J1_122_2300_n103 MAJIxp5_ASAP7_75t_R
XU287 VSS VDD  n192 n145 DP_OP_10J1_122_2300_n219 NOR2x1_ASAP7_75t_R
XU288 VSS VDD  DP_OP_10J1_122_2300_n101 DP_OP_10J1_122_2300_n98 DP_OP_10J1_122_2300_n79 n205 MAJIxp5_ASAP7_75t_R
XU289 VSS VDD  n187 n206 n188 NAND2xp5_ASAP7_75t_R
XU290 VSS VDD  n191 n190 n220 XOR2xp5_ASAP7_75t_R
XU291 VSS VDD  n129 n154 n219 NOR2xp33_ASAP7_75t_R
XU292 VSS VDD  n121 n219 n220 n224 MAJIxp5_ASAP7_75t_R
XU293 VSS VDD  n194 n193 n195 XOR2xp5_ASAP7_75t_R
XU294 VSS VDD  n196 n195 n222 XNOR2xp5_ASAP7_75t_R
XU295 VSS VDD  n198 n197 n200 XOR2xp5_ASAP7_75t_R
XU296 VSS VDD  n200 n199 n221 XNOR2xp5_ASAP7_75t_R
XU297 VSS VDD  n224 n222 n221 n226 MAJIxp5_ASAP7_75t_R
XU298 VSS VDD  DP_OP_10J1_122_2300_n120 DP_OP_10J1_122_2300_n140 DP_OP_10J1_122_2300_n122 n204 MAJIxp5_ASAP7_75t_R
XU299 VSS VDD  n133 n204 n202 XNOR2xp5_ASAP7_75t_R
XU300 VSS VDD  n205 DP_OP_10J1_122_2300_n53 n207 XNOR2xp5_ASAP7_75t_R
XU301 VSS VDD  In_Weight_4[0] In_IFM_4[3] n214 NAND2x1p5_ASAP7_75t_R
XU302 VSS VDD  In_Weight_4[0] In_IFM_4[2] DP_OP_10J1_122_2300_n175 AND2x4_ASAP7_75t_R
XU303 VSS VDD  n164 n243 DP_OP_10J1_122_2300_n192 NOR2xp33_ASAP7_75t_R
XU304 VSS VDD  n118 n183 DP_OP_10J1_122_2300_n216 NOR2xp33_ASAP7_75t_R
XU305 VSS VDD  In_Weight_3[0] n242 INVx8_ASAP7_75t_R
XU306 VSS VDD  n242 n124 DP_OP_10J1_122_2300_n243 NOR2xp33_ASAP7_75t_R
XU307 VSS VDD  n220 n219 n147 A5  Out_OFM[0] FAx1_ASAP7_75t_R
XU308 VSS VDD  n222 n221 n223 XOR2xp5_ASAP7_75t_R
XU309 VSS VDD  n224 n223 A6  Out_OFM[1] HAxp5_ASAP7_75t_R
XU310 VSS VDD  DP_OP_10J1_122_2300_n143 DP_OP_10J1_122_2300_n141 A7  n225 HAxp5_ASAP7_75t_R
XU311 VSS VDD  n226 n225 A8  Out_OFM[2] HAxp5_ASAP7_75t_R
XU312 VSS VDD  n230 n229 A9  Out_OFM[3] HAxp5_ASAP7_75t_R
XU313 VSS VDD  n233 n232 A10  DP_OP_10J1_122_2300_n51 HAxp5_ASAP7_75t_R
XU314 VSS VDD  In_IFM_4[3] In_Weight_4[2] n235 NAND2x1p5_ASAP7_75t_R
XU315 VSS VDD  n235 n234 A11  DP_OP_10J1_122_2300_n70 HAxp5_ASAP7_75t_R
XU316 VSS VDD  n238 n237 DP_OP_10J1_122_2300_n73 OR2x2_ASAP7_75t_R
XU317 VSS VDD  n235 n234 DP_OP_10J1_122_2300_n80 NOR2xp33_ASAP7_75t_R
XU318 VSS VDD  In_Weight_4[1] In_IFM_4[1] DP_OP_10J1_122_2300_n178 AND2x4_ASAP7_75t_R
XU319 VSS VDD  DP_OP_10J1_122_2300_n41 n150 n246 XOR2xp5_ASAP7_75t_R
XU320 VSS VDD  n210 n30 n247 XNOR2xp5_ASAP7_75t_R
XU321 VSS VDD  n107 DP_OP_10J1_122_2300_n64 A12  n249 HAxp5_ASAP7_75t_R
.ENDS


