.TITLE Comparator
*****************************
**     Library setting     **
*****************************
.protect
.include '7nm_TT.pm'
.include 'asap7sc7p5t_INVBUF_RVT.sp'
.include 'asap7sc7p5t_SIMPLE_RVT.sp'
.include 'Buffer.sp'
.unprotect
*.param   VDD_c = 0.4
.vec 'Pattern_convolution.vec'
*****************************
**     Voltage Source      **
*****************************
.global VDD GND
VDD VDD GND 0.4
xbuf0  IFM0_0 IFM0_0_ buffer
xbuf1  IFM0_1 IFM0_1_ buffer
xbuf2  IFM0_2 IFM0_2_ buffer
xbuf3  IFM0_3 IFM0_3_ buffer
xbuf4  IFM1_0 IFM1_0_ buffer
xbuf5  IFM1_1 IFM1_1_ buffer
xbuf6  IFM1_2 IFM1_2_ buffer
xbuf7  IFM1_3 IFM1_3_ buffer
xbuf8  IFM2_0 IFM2_0_ buffer
xbuf9  IFM2_1 IFM2_1_ buffer
xbuf10 IFM2_2 IFM2_2_ buffer
xbuf11 IFM2_3 IFM2_3_ buffer
xbuf12 IFM3_0 IFM3_0_ buffer
xbuf13 IFM3_1 IFM3_1_ buffer
xbuf14 IFM3_2 IFM3_2_ buffer
xbuf15 IFM3_3 IFM3_3_ buffer

xbuf16 INW0_0 INW0_0_ buffer
xbuf17 INW0_1 INW0_1_ buffer
xbuf18 INW0_2 INW0_2_ buffer
xbuf19 INW0_3 INW0_3_ buffer
xbuf20 INW1_0 INW1_0_ buffer
xbuf21 INW1_1 INW1_1_ buffer
xbuf22 INW1_2 INW1_2_ buffer
xbuf23 INW1_3 INW1_3_ buffer
xbuf24 INW2_0 INW2_0_ buffer
xbuf25 INW2_1 INW2_1_ buffer
xbuf26 INW2_2 INW2_2_ buffer
xbuf27 INW2_3 INW2_3_ buffer
xbuf28 INW3_0 INW3_0_ buffer
xbuf29 INW3_1 INW3_1_ buffer
xbuf30 INW3_2 INW3_2_ buffer
xbuf31 INW3_3 INW3_3_ buffer

cout0 out0 GND 5f
cout1 out1 GND 5f
cout2 out2 GND 5f
cout3 out3 GND 5f
cout4 out4 GND 5f
cout5 out5 GND 5f
cout6 out6 GND 5f
cout7 out7 GND 5f
cout8 out8 GND 5f
cout9 out9 GND 5f

xConvolution GND VDD IFM0_3_ IFM0_2_ IFM0_1_ IFM0_0_ IFM1_3_ IFM1_2_ IFM1_1_ IFM1_0_ IFM2_3_ IFM2_2_ IFM2_1_ IFM2_0_ IFM3_3_ IFM3_2_ IFM3_1_ IFM3_0_ INW0_3_ INW0_2_ INW0_1_ INW0_0_ INW1_3_ INW1_2_ INW1_1_ INW1_0_ INW2_3_ INW2_2_ INW2_1_ INW2_0_ INW3_3_ INW3_2_ INW3_1_ INW3_0_ out9 out8 out7 out6 out5 out4 out3 out2 out1 out0 Convolution
.SUBCKT Convolution VSS VDD  IFM_0[3] IFM_0[2] IFM_0[1] IFM_0[0] IFM_1[3] IFM_1[2] IFM_1[1] IFM_1[0] IFM_2[3] IFM_2[2] IFM_2[1] IFM_2[0] IFM_3[3] IFM_3[2] IFM_3[1] IFM_3[0] INW_0[3] INW_0[2] INW_0[1] INW_0[0] INW_1[3] INW_1[2] INW_1[1] INW_1[0] INW_2[3] INW_2[2] INW_2[1] INW_2[0] INW_3[3] INW_3[2] INW_3[1] INW_3[0] Output[9] Output[8] Output[7] Output[6] Output[5] Output[4] Output[3] Output[2] Output[1] Output[0]
Xmult_19 VSS VDD  IFM_0[3] IFM_0[2] IFM_0[1] IFM_0[0] INW_0[3] INW_0[2] INW_0[1] INW_0[0] N7 N6 N5 N4 N3 N2 N1 N0 Convolution_DW_mult_uns_3
Xmult_19_2 VSS VDD  IFM_1[3] IFM_1[2] IFM_1[1] IFM_1[0] INW_1[3] INW_1[2] INW_1[1] INW_1[0] N15 N14 N13 N12 N11 N10 N9 N8 Convolution_DW_mult_uns_2
Xmult_19_3 VSS VDD  IFM_2[3] IFM_2[2] IFM_2[1] IFM_2[0] INW_2[3] INW_2[2] INW_2[1] INW_2[0] N32 N31 N30 N29 N28 N27 N26 N25 Convolution_DW_mult_uns_1
Xmult_19_4 VSS VDD  IFM_3[3] IFM_3[2] IFM_3[1] IFM_3[0] INW_3[3] INW_3[2] INW_3[1] INW_3[0] N50 N49 N48 N47 N46 N45 N44 N43 Convolution_DW_mult_uns_0
Xadd_1_root_add_0_root_add_19_3 VSS VDD  N42 N42 N15 N14 N13 N12 N11 N10 N9 N8 N42 N42 N50 N49 N48 N47 N46 N45 N44 N43 N42 GND net9 net8 net7 net6 net5 net4 net3 net2 net1 Convolution_DW01_add_2
Xadd_2_root_add_0_root_add_19_3 VSS VDD  N42 N42 N7 N6 N5 N4 N3 N2 N1 N0 N42 N42 N32 N31 N30 N29 N28 N27 N26 N25 N42 GND N41 N40 N39 N38 N37 N36 N35 N34 N33 Convolution_DW01_add_1
Xadd_0_root_add_0_root_add_19_3 VSS VDD  N42 N41 N40 N39 N38 N37 N36 N35 N34 N33 N42 net9 net8 net7 net6 net5 net4 net3 net2 net1 N42 Output[9] Output[8] Output[7] Output[6] Output[5] Output[4] Output[3] Output[2] Output[1] Output[0] Convolution_DW01_add_0
XU1 VSS VDD  N42 TIELOx1_ASAP7_75t_R
.ENDS


.SUBCKT  Convolution_DW01_add_0 VSS VDD A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CI SUM[9] SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0] 
XU1_8 VSS VDD  A[8] B[8] n3 n10 n11 FAx1_ASAP7_75t_R
XU1_7 VSS VDD  A[7] B[7] n4 n12 n13 FAx1_ASAP7_75t_R
XU1_6 VSS VDD  A[6] B[6] n5 n14 n15 FAx1_ASAP7_75t_R
XU1_5 VSS VDD  A[5] B[5] n6 n16 n17 FAx1_ASAP7_75t_R
XU1_4 VSS VDD  A[4] B[4] n7 n18 n19 FAx1_ASAP7_75t_R
XU1_3 VSS VDD  A[3] B[3] n8 n20 n21 FAx1_ASAP7_75t_R
XU1_2 VSS VDD  A[2] B[2] n9 n22 n23 FAx1_ASAP7_75t_R
XU1_1 VSS VDD  A[1] B[1] n1 n24 n25 FAx1_ASAP7_75t_R
XU1 VSS VDD  A[0] B[0] n1 AND2x2_ASAP7_75t_R
XU2 VSS VDD  B[0] A[0] SUM[0] XOR2xp5_ASAP7_75t_R
XU3 VSS VDD  n12 n3 INVx1_ASAP7_75t_R
XU4 VSS VDD  n14 n4 INVx1_ASAP7_75t_R
XU5 VSS VDD  n16 n5 INVx1_ASAP7_75t_R
XU6 VSS VDD  n18 n6 INVx1_ASAP7_75t_R
XU7 VSS VDD  n20 n7 INVx1_ASAP7_75t_R
XU8 VSS VDD  n22 n8 INVx1_ASAP7_75t_R
XU9 VSS VDD  n24 n9 INVx1_ASAP7_75t_R
XU10 VSS VDD  n10 SUM[9] INVx1_ASAP7_75t_R
XU11 VSS VDD  n11 SUM[8] INVx1_ASAP7_75t_R
XU12 VSS VDD  n13 SUM[7] INVx1_ASAP7_75t_R
XU13 VSS VDD  n15 SUM[6] INVx1_ASAP7_75t_R
XU14 VSS VDD  n17 SUM[5] INVx1_ASAP7_75t_R
XU15 VSS VDD  n19 SUM[4] INVx1_ASAP7_75t_R
XU16 VSS VDD  n21 SUM[3] INVx1_ASAP7_75t_R
XU17 VSS VDD  n23 SUM[2] INVx1_ASAP7_75t_R
XU18 VSS VDD  n25 SUM[1] INVx1_ASAP7_75t_R
.ENDS


.SUBCKT   Convolution_DW01_add_1  VSS VDD A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CI SUM[9] SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0]
XU1_7 VSS VDD  A[7] B[7] n3 n9 n10 FAx1_ASAP7_75t_R
XU1_6 VSS VDD  A[6] B[6] n4 n11 n12 FAx1_ASAP7_75t_R
XU1_5 VSS VDD  A[5] B[5] n5 n13 n14 FAx1_ASAP7_75t_R
XU1_4 VSS VDD  A[4] B[4] n6 n15 n16 FAx1_ASAP7_75t_R
XU1_3 VSS VDD  A[3] B[3] n7 n17 n18 FAx1_ASAP7_75t_R
XU1_2 VSS VDD  A[2] B[2] n8 n19 n20 FAx1_ASAP7_75t_R
XU1_1 VSS VDD  A[1] B[1] n2 n21 n22 FAx1_ASAP7_75t_R
XU1 VSS VDD  B[0] A[0] SUM[0] XOR2xp5_ASAP7_75t_R
XU2 VSS VDD  A[0] B[0] n2 AND2x2_ASAP7_75t_R
XU3 VSS VDD  n11 n3 INVx1_ASAP7_75t_R
XU4 VSS VDD  n13 n4 INVx1_ASAP7_75t_R
XU5 VSS VDD  n15 n5 INVx1_ASAP7_75t_R
XU6 VSS VDD  n17 n6 INVx1_ASAP7_75t_R
XU7 VSS VDD  n19 n7 INVx1_ASAP7_75t_R
XU8 VSS VDD  n21 n8 INVx1_ASAP7_75t_R
XU9 VSS VDD  n9 SUM[8] INVx1_ASAP7_75t_R
XU10 VSS VDD  n10 SUM[7] INVx1_ASAP7_75t_R
XU11 VSS VDD  n12 SUM[6] INVx1_ASAP7_75t_R
XU12 VSS VDD  n14 SUM[5] INVx1_ASAP7_75t_R
XU13 VSS VDD  n16 SUM[4] INVx1_ASAP7_75t_R
XU14 VSS VDD  n18 SUM[3] INVx1_ASAP7_75t_R
XU15 VSS VDD  n20 SUM[2] INVx1_ASAP7_75t_R
XU16 VSS VDD  n22 SUM[1] INVx1_ASAP7_75t_R
.ENDS


.SUBCKT  Convolution_DW01_add_2 VSS VDD  A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CI SUM[9] SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0]
XU1_7 VSS VDD  A[7] B[7] n3 n9 n10 FAx1_ASAP7_75t_R
XU1_6 VSS VDD  A[6] B[6] n4 n11 n12 FAx1_ASAP7_75t_R
XU1_5 VSS VDD  A[5] B[5] n5 n13 n14 FAx1_ASAP7_75t_R
XU1_4 VSS VDD  A[4] B[4] n6 n15 n16 FAx1_ASAP7_75t_R
XU1_3 VSS VDD  A[3] B[3] n7 n17 n18 FAx1_ASAP7_75t_R
XU1_2 VSS VDD  A[2] B[2] n8 n19 n20 FAx1_ASAP7_75t_R
XU1_1 VSS VDD  A[1] B[1] n1 n21 n22 FAx1_ASAP7_75t_R
XU1 VSS VDD  A[0] B[0] n1 AND2x2_ASAP7_75t_R
XU2 VSS VDD  B[0] A[0] SUM[0] XOR2xp5_ASAP7_75t_R
XU3 VSS VDD  n11 n3 INVx1_ASAP7_75t_R
XU4 VSS VDD  n13 n4 INVx1_ASAP7_75t_R
XU5 VSS VDD  n15 n5 INVx1_ASAP7_75t_R
XU6 VSS VDD  n17 n6 INVx1_ASAP7_75t_R
XU7 VSS VDD  n19 n7 INVx1_ASAP7_75t_R
XU8 VSS VDD  n21 n8 INVx1_ASAP7_75t_R
XU9 VSS VDD  n9 SUM[8] INVx1_ASAP7_75t_R
XU10 VSS VDD  n10 SUM[7] INVx1_ASAP7_75t_R
XU11 VSS VDD  n12 SUM[6] INVx1_ASAP7_75t_R
XU12 VSS VDD  n14 SUM[5] INVx1_ASAP7_75t_R
XU13 VSS VDD  n16 SUM[4] INVx1_ASAP7_75t_R
XU14 VSS VDD  n18 SUM[3] INVx1_ASAP7_75t_R
XU15 VSS VDD  n20 SUM[2] INVx1_ASAP7_75t_R
XU16 VSS VDD  n22 SUM[1] INVx1_ASAP7_75t_R
.ENDS


.SUBCKT   Convolution_DW_mult_uns_0 VSS VDD a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 VSS VDD  n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 VSS VDD  n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 VSS VDD  n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 VSS VDD  a[2] n83 INVx1_ASAP7_75t_R
XU71 VSS VDD  n35 n84 INVx1_ASAP7_75t_R
XU72 VSS VDD  a[0] n85 INVx1_ASAP7_75t_R
XU73 VSS VDD  b[3] n86 INVx1_ASAP7_75t_R
XU74 VSS VDD  b[0] n87 INVx1_ASAP7_75t_R
XU75 VSS VDD  n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 VSS VDD  n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 VSS VDD  n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 VSS VDD  n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 VSS VDD  n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 VSS VDD  b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 VSS VDD  n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 VSS VDD  n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 VSS VDD  n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 VSS VDD  n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 VSS VDD  n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 VSS VDD  n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 VSS VDD  n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 VSS VDD  n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 VSS VDD  n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 VSS VDD  n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 VSS VDD  n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 VSS VDD  n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 VSS VDD  n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 VSS VDD  n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 VSS VDD  n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 VSS VDD  n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 VSS VDD  n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 VSS VDD  n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 VSS VDD  n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 VSS VDD  n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 VSS VDD  n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 VSS VDD  n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 VSS VDD  n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 VSS VDD  n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 VSS VDD  n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 VSS VDD  b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 VSS VDD  b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 VSS VDD  n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 VSS VDD  n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 VSS VDD  a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 VSS VDD  a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 VSS VDD  n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 VSS VDD  b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 VSS VDD  n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 VSS VDD  b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 VSS VDD  b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 VSS VDD  n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 VSS VDD  a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 VSS VDD  a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 VSS VDD  n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 VSS VDD  n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 VSS VDD  a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 VSS VDD  b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT  Convolution_DW_mult_uns_1 VSS VDD  a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 VSS VDD  n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 VSS VDD  n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 VSS VDD  n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 VSS VDD  a[2] n83 INVx1_ASAP7_75t_R
XU71 VSS VDD  n35 n84 INVx1_ASAP7_75t_R
XU72 VSS VDD  a[0] n85 INVx1_ASAP7_75t_R
XU73 VSS VDD  b[3] n86 INVx1_ASAP7_75t_R
XU74 VSS VDD  b[0] n87 INVx1_ASAP7_75t_R
XU75 VSS VDD  n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 VSS VDD  n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 VSS VDD  n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 VSS VDD  n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 VSS VDD  n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 VSS VDD  b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 VSS VDD  n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 VSS VDD  n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 VSS VDD  n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 VSS VDD  n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 VSS VDD  n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 VSS VDD  n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 VSS VDD  n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 VSS VDD  n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 VSS VDD  n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 VSS VDD  n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 VSS VDD  n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 VSS VDD  n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 VSS VDD  n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 VSS VDD  n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 VSS VDD  n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 VSS VDD  n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 VSS VDD  n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 VSS VDD  n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 VSS VDD  n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 VSS VDD  n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 VSS VDD  n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 VSS VDD  n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 VSS VDD  n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 VSS VDD  n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 VSS VDD  n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 VSS VDD  b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 VSS VDD  b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 VSS VDD  n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 VSS VDD  n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 VSS VDD  a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 VSS VDD  a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 VSS VDD  n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 VSS VDD  b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 VSS VDD  n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 VSS VDD  b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 VSS VDD  b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 VSS VDD  n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 VSS VDD  a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 VSS VDD  a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 VSS VDD  n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 VSS VDD  n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 VSS VDD  a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 VSS VDD  b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT   Convolution_DW_mult_uns_2 VSS VDD a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 VSS VDD  n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 VSS VDD  n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 VSS VDD  n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 VSS VDD  a[2] n83 INVx1_ASAP7_75t_R
XU71 VSS VDD  n35 n84 INVx1_ASAP7_75t_R
XU72 VSS VDD  a[0] n85 INVx1_ASAP7_75t_R
XU73 VSS VDD  b[3] n86 INVx1_ASAP7_75t_R
XU74 VSS VDD  b[0] n87 INVx1_ASAP7_75t_R
XU75 VSS VDD  n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 VSS VDD  n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 VSS VDD  n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 VSS VDD  n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 VSS VDD  n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 VSS VDD  b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 VSS VDD  n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 VSS VDD  n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 VSS VDD  n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 VSS VDD  n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 VSS VDD  n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 VSS VDD  n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 VSS VDD  n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 VSS VDD  n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 VSS VDD  n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 VSS VDD  n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 VSS VDD  n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 VSS VDD  n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 VSS VDD  n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 VSS VDD  n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 VSS VDD  n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 VSS VDD  n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 VSS VDD  n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 VSS VDD  n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 VSS VDD  n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 VSS VDD  n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 VSS VDD  n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 VSS VDD  n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 VSS VDD  n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 VSS VDD  n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 VSS VDD  n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 VSS VDD  b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 VSS VDD  b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 VSS VDD  n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 VSS VDD  n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 VSS VDD  a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 VSS VDD  a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 VSS VDD  n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 VSS VDD  b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 VSS VDD  n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 VSS VDD  b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 VSS VDD  b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 VSS VDD  n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 VSS VDD  a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 VSS VDD  a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 VSS VDD  n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 VSS VDD  n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 VSS VDD  a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 VSS VDD  b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT  Convolution_DW_mult_uns_3  VSS VDD a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 VSS VDD  n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 VSS VDD  n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 VSS VDD  n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 VSS VDD  a[2] n83 INVx1_ASAP7_75t_R
XU71 VSS VDD  n35 n84 INVx1_ASAP7_75t_R
XU72 VSS VDD  a[0] n85 INVx1_ASAP7_75t_R
XU73 VSS VDD  b[3] n86 INVx1_ASAP7_75t_R
XU74 VSS VDD  b[0] n87 INVx1_ASAP7_75t_R
XU75 VSS VDD  n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 VSS VDD  n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 VSS VDD  n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 VSS VDD  n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 VSS VDD  n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 VSS VDD  b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 VSS VDD  n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 VSS VDD  n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 VSS VDD  n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 VSS VDD  n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 VSS VDD  n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 VSS VDD  n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 VSS VDD  n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 VSS VDD  n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 VSS VDD  n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 VSS VDD  n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 VSS VDD  n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 VSS VDD  n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 VSS VDD  n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 VSS VDD  n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 VSS VDD  n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 VSS VDD  n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 VSS VDD  n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 VSS VDD  n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 VSS VDD  n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 VSS VDD  n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 VSS VDD  n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 VSS VDD  n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 VSS VDD  n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 VSS VDD  n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 VSS VDD  n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 VSS VDD  b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 VSS VDD  b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 VSS VDD  n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 VSS VDD  n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 VSS VDD  a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 VSS VDD  a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 VSS VDD  n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 VSS VDD  b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 VSS VDD  n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 VSS VDD  b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 VSS VDD  b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 VSS VDD  n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 VSS VDD  a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 VSS VDD  a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 VSS VDD  n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 VSS VDD  n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 VSS VDD  a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 VSS VDD  b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS



*****************************
**      Measurement        **
*****************************
.tran 0.01ns 100ns 0.01ns
.measure TRAN delay  TRIG V(INW3_2_) VAL=0.2 FALL=1 TARG V(out8) VAL=0.2 RISE=2
* .measure TRAN TR     TRIG V(out) VAL=0.04 RISE=1 TARG V(out) VAL=0.36 RISE=1
* .measure TRAN TF     TRIG V(out) VAL=0.36 FALL=1 TARG V(out) VAL=0.04 FALL=1
.meas tran pwr avg POWER 

*** 
*****************************
**    Simulator setting    **
*****************************
.option post 
.options probe	
.probe v(INW*_) v(IFM*_) v(out*)
.option captab	
.TEMP 25

.op

.end